// prosys.v

// Generated using ACDS version 16.1 196

`timescale 1 ps / 1 ps
module prosys (
		input  wire  clk_clk,       //   clk.clk
		input  wire  reset_reset_n  // reset.reset_n
	);

endmodule
